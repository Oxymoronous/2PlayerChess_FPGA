module mouse_rom ( input [3:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 4;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		16'b1110000000000000,
		16'b1111100000000000,
		16'b1111110000000000,
		16'b1111111100000000,
		16'b1111111110000000,
		16'b1111111111000000,
		16'b1111111111100000,
		16'b1111111111110000,
		16'b1111111111111000,
		16'b1111111111111100,
		16'b1111111111111110,
		16'b1111111111111111,
		16'b1111111111000000,
		16'b1110001111100000,
		16'b1100000111110000,
		16'b0000000011111000
	};
	
	assign data = ROM[addr];
	
endmodule
